`timescale 1ns/1ps

module testbench;

    reg [63:0] a;
    reg [63:0] b;

    wire [63:0] s;

    barrel_shifter_left uut (.data(a), ._shift(b), .out(s));

    initial begin
    
        $dumpfile("GTK/barrel_left64bit.vcd");
        $dumpvars(0, testbench);

        // Gpt generated test cases - 


        a = 64'h0000_0000_0000_0001;

        // -------------------------
        // Test 1: shift = 0
        // -------------------------
        b = 64'd0;
        #10;

        // -------------------------
        // Test 2: shift = 1
        // -------------------------
        b = 64'd1;
        #10;

        // -------------------------
        // Test 3: shift = 4
        // -------------------------
        b = 64'd4;
        #10;

        // -------------------------
        // Test 4: shift = 13 (8+4+1)
        // -------------------------
        b = 64'd13;
        #10;

        // -------------------------
        // Test 5: shift = 32
        // -------------------------
        b = 64'd32;
        #10;

        // -------------------------
        // Test 6: shift = 63 (max)
        // -------------------------
        b = 64'd63;
        #10;

        // -------------------------
        // Test 6: shift = 65 (mask check)
        // -------------------------
        b = 64'd65;
        #10;


        // -------------------------
        // Test 9: complex pattern
        // -------------------------
        a = 64'hF0F0_F0F0_F0F0_F0F0;
        b = 64'd4;
        #10;

        // -------------------------
        // Test 10: MSB test
        // -------------------------
        a = 64'h8000_0000_0000_0000;
        b = 64'd1;
        #10;

        $finish;
     
    end

endmodule