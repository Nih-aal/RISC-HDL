`timescale 1ns/1ps

module testbench;

    reg [63:0] a;
    reg [63:0] b;

    wire [63:0] s;

    barrel_shifter_right_logical uut (.data(a), ._shift(b), .out(s));

    initial begin
    
        $dumpfile("GTK/barrel_logical_right64bit.vcd");
        $dumpvars(0, testbench);

        // Gpt generated test cases - 

        a = 64'h8000000000000000;

        // --------------------------------
        // Test 1: shift = 0 (identity)
        // --------------------------------
        
        b = 64'd0;
        #10;

        // --------------------------------
        // Test 2: shift = 1
        // --------------------------------
        b = 64'd1;
        #10;

        // --------------------------------
        // Test 3: shift = 4
        // --------------------------------
        b = 64'd4;
        #10;

        // --------------------------------
        // Test 4: shift = 13 (8+4+1)
        // --------------------------------
        b = 64'd13;
        #10;

        // --------------------------------
        // Test 5: shift = 32
        // --------------------------------
        b = 64'd32;
        #10;

        // --------------------------------
        // Test 6: shift = 63 (max)
        // --------------------------------
        b = 64'd63;
        #10;

        // --------------------------------
        // Test 7: shift = 65 (mask check)
        // --------------------------------
        b = 64'd65;
        #10;

        // --------------------------------
        // Test 8: single-bit LSB pattern
        // --------------------------------
        a = 64'h0000_0000_0000_0001;
        b = 64'd1;
        #10;

        // --------------------------------
        // Test 10: alternating pattern
        // --------------------------------
        a = 64'hA0A0_A0A0_A0A0_A0A0;
        b = 64'd4;
        #10;

        $finish;
     
    end

endmodule